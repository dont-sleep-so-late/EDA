LIBRARY IEEE;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY encode_BCD IS
PORT(
	hexin :IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	BCDOUT: OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
	);
END encode_BCD;

ARCHITECTURE RTL OF encode_BCD IS
BEGIN
	PROCESS(hexin)
	VARIABLE NUM :INTEGER RANGE 0 TO 255;
	VARIABLE HUNDRED,TEN,ONE :INTEGER RANGE 0 TO 9;
	VARIABLE H,T,O :STD_LOGIC_VECTOR(3 DOWNTO 0);
	BEGIN
	NUM:=CONV_INTEGER(hexin);
	HUNDRED:=NUM/100;
	TEN:=(NUM MOD 100)/10;
	ONE:=NUM MOD 10;
	H:=CONV_STD_LOGIC_VECTOR(HUNDRED,4);
	T:=CONV_STD_LOGIC_VECTOR(TEN,4);
	O:=CONV_STD_LOGIC_VECTOR(ONE,4);
	BCDOUT<=H&T&O;
	END PROCESS;
END RTL;